`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/12/01 15:24:56
// Design Name: 
// Module Name: pipeline_md5
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pipeline_md5(
    input clk,
    //input st,
    input [63:0] num,
    //input [127:0] hash,
    output reg[127:0] answer,
    output reg [63:0] currnum
    //output done
    );
reg [31:0] a,a0, a1, a2, a3, a4, a5, a6, a7, a8, a9,a10,a11,a12,a13,a14,a15,a16,
              a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31,a32,
              a33,a34,a35,a36,a37,a38,a39,a40,a41,a42,a43,a44,a45,a46,a47,a48,
              a49,a50,a51,a52,a53,a54,a55,a56,a57,a58,a59,a60,a61,a62,a63,a64 = 0;
reg [31:0] b,b0, b1, b2, b3, b4, b5, b6, b7, b8, b9,b10,b11,b12,b13,b14,b15,b16,
              b17,b18,b19,b20,b21,b22,b23,b24,b25,b26,b27,b28,b29,b30,b31,b32,
              b33,b34,b35,b36,b37,b38,b39,b40,b41,b42,b43,b44,b45,b46,b47,b48,
              b49,b50,b51,b52,b53,b54,b55,b56,b57,b58,b59,b60,b61,b62,b63,b64 = 0;
reg [31:0] c,c0, c1, c2, c3, c4, c5, c6, c7, c8, c9,c10,c11,c12,c13,c14,c15,c16,
              c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,c31,c32,
              c33,c34,c35,c36,c37,c38,c39,c40,c41,c42,c43,c44,c45,c46,c47,c48,
              c49,c50,c51,c52,c53,c54,c55,c56,c57,c58,c59,c60,c61,c62,c63,c64 = 0;
reg [31:0] d,d0, d1, d2, d3, d4, d5, d6, d7, d8, d9,d10,d11,d12,d13,d14,d15,d16,
              d17,d18,d19,d20,d21,d22,d23,d24,d25,d26,d27,d28,d29,d30,d31,d32,
              d33,d34,d35,d36,d37,d38,d39,d40,d41,d42,d43,d44,d45,d46,d47,d48,
              d49,d50,d51,d52,d53,d54,d55,d56,d57,d58,d59,d60,d61,d62,d63,d64 = 0;
reg [63:0] n,n0, n1, n2, n3, n4, n5, n6, n7, n8, n9,n10,n11,n12,n13,n14,n15,n16,
              n17,n18,n19,n20,n21,n22,n23,n24,n25,n26,n27,n28,n29,n30,n31,n32,
              n33,n34,n35,n36,n37,n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,
              n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64 = 0;
reg [31:0] e0 = 32'h00000080;        
reg [31:0] e1 = 32'h00000040;

//assign answer = {a64[7:0],a64[15:8],a64[23:16],a64[31:24],
//                 b64[7:0],b64[15:8],b64[23:16],b64[31:24],
//                 c64[7:0],c64[15:8],c64[23:16],c64[31:24],
//                 d64[7:0],d64[15:8],d64[23:16],d64[31:24]};
//assign currnum = {n64[39:32],n64[47:40],n64[55:48],n64[63:56],
//                  n64[7:0],n64[15:8],n64[23:16],n64[31:24]};

always@(posedge clk) begin 
        answer <= {a64[7:0],a64[15:8],a64[23:16],a64[31:24],
                 b64[7:0],b64[15:8],b64[23:16],b64[31:24],
                 c64[7:0],c64[15:8],c64[23:16],c64[31:24],
                 d64[7:0],d64[15:8],d64[23:16],d64[31:24]};
        currnum <= {n64[39:32],n64[47:40],n64[55:48],n64[63:56],
                  n64[7:0],n64[15:8],n64[23:16],n64[31:24]};
        a <= 32'h67452301;
        b <= 32'hefcdab89;
        c <= 32'h98badcfe;
        d <= 32'h10325476;
        //n <= "43218765";
        //num "12345678"
        n <= {num[39:32],num[47:40],num[55:48],num[63:56],
              num[7:0],num[15:8],num[23:16],num[31:24]};
        

        a10 <= d9; a9 <= d8; a8 <= d7; a7 <= d6; a6 <= d5; a5 <= d4; a4 <= d3; a3 <= d2; a2 <= d1; a1 <= d0; a0 <= d;
        a20 <= d19; a19 <= d18; a18 <= d17; a17 <= d16; a16 <= d15; a15 <= d14; a14 <= d13; a13 <= d12; a12 <= d11; a11 <= d10;
        a30 <= d29; a29 <= d28; a28 <= d27; a27 <= d26; a26 <= d25; a25 <= d24; a24 <= d23; a23 <= d22; a22 <= d21; a21 <= d20;
        a40 <= d39; a39 <= d38; a38 <= d37; a37 <= d36; a36 <= d35; a35 <= d34; a34 <= d33; a33 <= d32; a32 <= d31; a31 <= d30;
        a50 <= d49; a49 <= d48; a48 <= d47; a47 <= d46; a46 <= d45; a45 <= d44; a44 <= d43; a43 <= d42; a42 <= d41; a41 <= d40;
        a60 <= d59; a59 <= d58; a58 <= d57; a57 <= d56; a56 <= d55; a55 <= d54; a54 <= d53; a53 <= d52; a52 <= d51; a51 <= d50;
        a63 <= d62; a62 <= d61; a61 <= d60;
        
        c10 <= b9; c9 <= b8; c8 <= b7; c7 <= b6; c6 <= b5; c5 <= b4; c4 <= b3; c3 <= b2; c2 <= b1; c1 <= b0; c0 <= b;
        c20 <= b19; c19 <= b18; c18 <= b17; c17 <= b16; c16 <= b15; c15 <= b14; c14 <= b13; c13 <= b12; c12 <= b11; c11 <= b10;
        c30 <= b29; c29 <= b28; c28 <= b27; c27 <= b26; c26 <= b25; c25 <= b24; c24 <= b23; c23 <= b22; c22 <= b21; c21 <= b20;
        c40 <= b39; c39 <= b38; c38 <= b37; c37 <= b36; c36 <= b35; c35 <= b34; c34 <= b33; c33 <= b32; c32 <= b31; c31 <= b30;
        c50 <= b49; c49 <= b48; c48 <= b47; c47 <= b46; c46 <= b45; c45 <= b44; c44 <= b43; c43 <= b42; c42 <= b41; c41 <= b40;
        c60 <= b59; c59 <= b58; c58 <= b57; c57 <= b56; c56 <= b55; c55 <= b54; c54 <= b53; c53 <= b52; c52 <= b51; c51 <= b50;
        c63 <= b62; c62 <= b61; c61 <= b60;
        
        d10 <= c9; d9 <= c8; d8 <= c7; d7 <= c6; d6 <= c5; d5 <= c4; d4 <= c3; d3 <= c2; d2 <= c1; d1 <= c0; d0 <= c;
        d20 <= c19; d19 <= c18; d18 <= c17; d17 <= c16; d16 <= c15; d15 <= c14; d14 <= c13; d13 <= c12; d12 <= c11; d11 <= c10;
        d30 <= c29; d29 <= c28; d28 <= c27; d27 <= c26; d26 <= c25; d25 <= c24; d24 <= c23; d23 <= c22; d22 <= c21; d21 <= c20;
        d40 <= c39; d39 <= c38; d38 <= c37; d37 <= c36; d36 <= c35; d35 <= c34; d34 <= c33; d33 <= c32; d32 <= c31; d31 <= c30;
        d50 <= c49; d49 <= c48; d48 <= c47; d47 <= c46; d46 <= c45; d45 <= c44; d44 <= c43; d43 <= c42; d42 <= c41; d41 <= c40;
        d60 <= c59; d59 <= c58; d58 <= c57; d57 <= c56; d56 <= c55; d55 <= c54; d54 <= c53; d53 <= c52; d52 <= c51; d51 <= c50;
        d63 <= c62; d62 <= c61; d61 <= c60;
        n0 <= n;
        n1 <= n0; n2 <= n1; n3 <= n2; n4 <= n3;
        n5 <= n4; n6 <= n5; n7 <= n6; n8 <= n7;
        n9 <= n8; n10 <= n9; n11 <= n10; n12 <= n11;
        n13 <= n12; n14 <= n13; n15 <= n14; n16 <= n15;
        n17 <= n16; n18 <= n17; n19 <= n18; n20 <= n19;
        n30 <= n29; n29 <= n28; n28 <= n27; n27 <= n26; n26 <= n25; n25 <= n24; n24 <= n23; n23 <= n22; n22 <= n21; n21 <= n20;
        n40 <= n39; n39 <= n38; n38 <= n37; n37 <= n36; n36 <= n35; n35 <= n34; n34 <= n33; n33 <= n32; n32 <= n31; n31 <= n30;
        n50 <= n49; n49 <= n48; n48 <= n47; n47 <= n46; n46 <= n45; n45 <= n44; n44 <= n43; n43 <= n42; n42 <= n41; n41 <= n40;
        n60 <= n59; n59 <= n58; n58 <= n57; n57 <= n56; n56 <= n55; n55 <= n54; n54 <= n53; n53 <= n52; n52 <= n51; n51 <= n50;
        n63 <= n62; n62 <= n61; n61 <= n60;
        n64 <= n63;
        //x = (a + ((b&c) | ((~b)&d)) + 32'hd76aa478 + n[31:0])
        b0 <= b + ((((a + ((b&c) | ((~b)&d)) + 32'hd76aa478 + n[63:32])) << 7) | (((a + ((b&c) | ((~b)&d)) + 32'hd76aa478 + n[63:32])) >> 32 - 7));
        b1 <= b0 + ((((a0 + ((b0&c0) | ((~b0)&d0)) + 32'he8c7b756 + n0[31:0])) << 12) | (((a0 + ((b0&c0) | ((~b0)&d0)) + 32'he8c7b756 + n0[31:0])) >> 32 - 12));
        b2 <= b1 + ((((a1 + ((b1&c1) | ((~b1)&d1)) + 32'h242070db + e0)) << 17) | (((a1 + ((b1&c1) | ((~b1)&d1)) + 32'h242070db + e0)) >> 32 - 17));
        b3 <= b2 + ((((a2 + ((b2&c2) | ((~b2)&d2)) + 32'hc1bdceee + 0)) << 22) | (((a2 + ((b2&c2) | ((~b2)&d2)) + 32'hc1bdceee + 0)) >> 32 - 22));
        
        b4 <= b3 + ((((a3 + ((b3&c3) | ((~b3)&d3)) + 32'hf57c0faf + 0)) << 7) | (((a3 + ((b3&c3) | ((~b3)&d3)) + 32'hf57c0faf + 0)) >> 32 - 7));
        b5 <= b4 + ((((a4 + ((b4&c4) | ((~b4)&d4)) + 32'h4787c62a + 0)) << 12) | (((a4 + ((b4&c4) | ((~b4)&d4)) + 32'h4787c62a + 0)) >> 32 - 12));
        b6 <= b5 + ((((a5 + ((b5&c5) | ((~b5)&d5)) + 32'ha8304613 + 0)) << 17) | (((a5 + ((b5&c5) | ((~b5)&d5)) + 32'ha8304613 + 0)) >> 32 - 17));
        b7 <= b6 + ((((a6 + ((b6&c6) | ((~b6)&d6)) + 32'hfd469501 + 0)) << 22) | (((a6 + ((b6&c6) | ((~b6)&d6)) + 32'hfd469501 + 0)) >> 32 - 22));
        
        b8 <= b7 + ((((a7 + ((b7&c7) | ((~b7)&d7)) + 32'h698098d8 + 0)) << 7) | (((a7 + ((b7&c7) | ((~b7)&d7)) + 32'h698098d8 + 0)) >> 32 - 7));
        b9 <= b8 + ((((a8 + ((b8&c8) | ((~b8)&d8)) + 32'h8b44f7af + 0)) << 12) | (((a8 + ((b8&c8) | ((~b8)&d8)) + 32'h8b44f7af + 0)) >> 32 - 12));
        b10 <= b9 + ((((a9 + ((b9&c9) | ((~b9)&d9)) + 32'hffff5bb1 + 0)) << 17) | (((a9 + ((b9&c9) | ((~b9)&d9)) + 32'hffff5bb1 + 0)) >> 32 - 17));
        b11 <= b10 + ((((a10 + ((b10&c10) | ((~b10)&d10)) + 32'h895cd7be + 0)) << 22) | (((a10 + ((b10&c10) | ((~b10)&d10)) + 32'h895cd7be + 0)) >> 32 - 22));
        
        b12 <= b11 + ((((a11 + ((b11&c11) | ((~b11)&d11)) + 32'h6b901122 + 0)) << 7) | (((a11 + ((b11&c11) | ((~b11)&d11)) + 32'h6b901122 + 0)) >> 32 - 7));
        b13 <= b12 + ((((a12 + ((b12&c12) | ((~b12)&d12)) + 32'hfd987193 + 0)) << 12) | (((a12 + ((b12&c12) | ((~b12)&d12)) + 32'hfd987193 + 0)) >> 32 - 12));
        b14 <= b13 + ((((a13 + ((b13&c13) | ((~b13)&d13)) + 32'ha679438e + e1)) << 17) | (((a13 + ((b13&c13) | ((~b13)&d13)) + 32'ha679438e + e1)) >> 32 - 17));
        b15 <= b14 + ((((a14 + ((b14&c14) | ((~b14)&d14)) + 32'h49b40821 + 0)) << 22) | (((a14 + ((b14&c14) | ((~b14)&d14)) + 32'h49b40821 + 0)) >> 32 - 22));
        
        //f = (d & b) | ((~d) & c);
        //g = (5*i + 1) % 16;
        b16 <= b15 + ((((a15 + ((d15 & b15) | ((~d15) & c15)) + 32'hf61e2562 + n15[31:0])) << 5) | (((a15 + ((d15 & b15) | ((~d15) & c15)) + 32'hf61e2562 + n15[31:0])) >> 32 - 5)); //g[1]
        b17 <= b16 + ((((a16 + ((d16 & b16) | ((~d16) & c16)) + 32'hc040b340 + 0)) << 9) | (((a16 + ((d16 & b16) | ((~d16) & c16)) + 32'hc040b340 + 0)) >> 32 - 9));
        b18 <= b17 + ((((a17 + ((d17 & b17) | ((~d17) & c17)) + 32'h265e5a51 + 0)) << 14) | (((a17 + ((d17 & b17) | ((~d17) & c17)) + 32'h265e5a51 + 0)) >> 32 - 14));
        b19 <= b18 + ((((a18 + ((d18 & b18) | ((~d18) & c18)) + 32'he9b6c7aa + n18[63:32])) << 20) | (((a18 + ((d18 & b18) | ((~d18) & c18)) + 32'he9b6c7aa + n18[63:32])) >> 32 - 20)); //g[0]
        
        b20 <= b19 + ((((a19 + ((d19 & b19) | ((~d19) & c19)) + 32'hd62f105d + 0)) << 5) | (((a19 + ((d19 & b19) | ((~d19) & c19)) + 32'hd62f105d + 0)) >> 32 - 5));
        b21 <= b20 + ((((a20 + ((d20 & b20) | ((~d20) & c20)) + 32'h02441453 + 0)) << 9) | (((a20 + ((d20 & b20) | ((~d20) & c20)) + 32'h02441453 + 0)) >> 32 - 9));
        b22 <= b21 + ((((a21 + ((d21 & b21) | ((~d21) & c21)) + 32'hd8a1e681 + 0)) << 14) | (((a21 + ((d21 & b21) | ((~d21) & c21)) + 32'hd8a1e681 + 0)) >> 32 - 14));
        b23 <= b22 + ((((a22 + ((d22 & b22) | ((~d22) & c22)) + 32'he7d3fbc8 + 0)) << 20) | (((a22 + ((d22 & b22) | ((~d22) & c22)) + 32'he7d3fbc8 + 0)) >> 32 - 20));
        
        b24 <= b23 + ((((a23 + ((d23 & b23) | ((~d23) & c23)) + 32'h21e1cde6 + 0)) << 5) | (((a23 + ((d23 & b23) | ((~d23) & c23)) + 32'h21e1cde6 + 0)) >> 32 - 5));
        b25 <= b24 + ((((a24 + ((d24 & b24) | ((~d24) & c24)) + 32'hc33707d6 + e1)) << 9) | (((a24 + ((d24 & b24) | ((~d24) & c24)) + 32'hc33707d6 + e1)) >> 32 - 9));
        b26 <= b25 + ((((a25 + ((d25 & b25) | ((~d25) & c25)) + 32'hf4d50d87 + 0)) << 14) | (((a25 + ((d25 & b25) | ((~d25) & c25)) + 32'hf4d50d87 + 0)) >> 32 - 14));
        b27 <= b26 + ((((a26 + ((d26 & b26) | ((~d26) & c26)) + 32'h455a14ed + 0)) << 20) | (((a26 + ((d26 & b26) | ((~d26) & c26)) + 32'h455a14ed + 0)) >> 32 - 20));
        
        b28 <= b27 + ((((a27 + ((d27 & b27) | ((~d27) & c27)) + 32'ha9e3e905 + 0)) << 5) | (((a27 + ((d27 & b27) | ((~d27) & c27)) + 32'ha9e3e905 + 0)) >> 32 - 5));
        b29 <= b28 + ((((a28 + ((d28 & b28) | ((~d28) & c28)) + 32'hfcefa3f8 + e0)) << 9) | (((a28 + ((d28 & b28) | ((~d28) & c28)) + 32'hfcefa3f8 + e0)) >> 32 - 9));
        b30 <= b29 + ((((a29 + ((d29 & b29) | ((~d29) & c29)) + 32'h676f02d9 + 0)) << 14) | (((a29 + ((d29 & b29) | ((~d29) & c29)) + 32'h676f02d9 + 0)) >> 32 - 14));
        b31 <= b30 + ((((a30 + ((d30 & b30) | ((~d30) & c30)) + 32'h8d2a4c8a + 0)) << 20) | (((a30 + ((d30 & b30) | ((~d30) & c30)) + 32'h8d2a4c8a + 0)) >> 32 - 20));
        
        //f = b ^ c ^ d;
        //g = (3*i + 5) % 16;
        b32 <= b31 + ((((a31 + (b31 ^ c31 ^ d31) + 32'hfffa3942 + 0)) << 4) | (((a31 + (b31 ^ c31 ^ d31) + 32'hfffa3942 + 0)) >> 32 - 4)); //
        b33 <= b32 + ((((a32 + (b32 ^ c32 ^ d32) + 32'h8771f681 + 0)) << 11) | (((a32 + (b32 ^ c32 ^ d32) + 32'h8771f681 + 0)) >> 32 - 11));
        b34 <= b33 + ((((a33 + (b33 ^ c33 ^ d33) + 32'h6d9d6122 + 0)) << 16) | (((a33 + (b33 ^ c33 ^ d33) + 32'h6d9d6122 + 0)) >> 32 - 16));
        b35 <= b34 + ((((a34 + (b34 ^ c34 ^ d34) + 32'hfde5380c + e1)) << 23) | (((a34 + (b34 ^ c34 ^ d34) + 32'hfde5380c + e1)) >> 32 - 23));
        
        b36 <= b35 + ((((a35 + (b35 ^ c35 ^ d35) + 32'ha4beea44 + n35[31:0])) << 4) | (((a35 + (b35 ^ c35 ^ d35) + 32'ha4beea44 + n35[31:0])) >> 32 - 4));  //g[1]
        b37 <= b36 + ((((a36 + (b36 ^ c36 ^ d36) + 32'h4bdecfa9 + 0)) << 11) | (((a36 + (b36 ^ c36 ^ d36) + 32'h4bdecfa9 + 0)) >> 32 - 11));
        b38 <= b37 + ((((a37 + (b37 ^ c37 ^ d37) + 32'hf6bb4b60 + 0)) << 16) | (((a37 + (b37 ^ c37 ^ d37) + 32'hf6bb4b60 + 0)) >> 32 - 16));
        b39 <= b38 + ((((a38 + (b38 ^ c38 ^ d38) + 32'hbebfbc70 + 0)) << 23) | (((a38 + (b38 ^ c38 ^ d38) + 32'hbebfbc70 + 0)) >> 32 - 23));
        
        b40 <= b39 + ((((a39 + (b39 ^ c39 ^ d39) + 32'h289b7ec6 + 0)) << 4) | (((a39 + (b39 ^ c39 ^ d39) + 32'h289b7ec6 + 0)) >> 32 - 4));
        b41 <= b40 + ((((a40 + (b40 ^ c40 ^ d40) + 32'heaa127fa + n40[63:32])) << 11) | (((a40 + (b40 ^ c40 ^ d40) + 32'heaa127fa + n40[63:32])) >> 32 - 11)); //g[0]
        b42 <= b41 + ((((a41 + (b41 ^ c41 ^ d41) + 32'hd4ef3085 + 0)) << 16) | (((a41 + (b41 ^ c41 ^ d41) + 32'hd4ef3085 + 0)) >> 32 - 16));
        b43 <= b42 + ((((a42 + (b42 ^ c42 ^ d42) + 32'h04881d05 + 0)) << 23) | (((a42 + (b42 ^ c42 ^ d42) + 32'h04881d05 + 0)) >> 32 - 23));
        
        b44 <= b43 + ((((a43 + (b43 ^ c43 ^ d43) + 32'hd9d4d039 + 0)) << 4) | (((a43 + (b43 ^ c43 ^ d43) + 32'hd9d4d039 + 0)) >> 32 - 4));
        b45 <= b44 + ((((a44 + (b44 ^ c44 ^ d44) + 32'he6db99e5 + 0)) << 11) | (((a44 + (b44 ^ c44 ^ d44) + 32'he6db99e5 + 0)) >> 32 - 11)); 
        b46 <= b45 + ((((a45 + (b45 ^ c45 ^ d45) + 32'h1fa27cf8 + 0)) << 16) | (((a45 + (b45 ^ c45 ^ d45) + 32'h1fa27cf8 + 0)) >> 32 - 16));
        b47 <= b46 + ((((a46 + (b46 ^ c46 ^ d46) + 32'hc4ac5665 + e0)) << 23) | (((a46 + (b46 ^ c46 ^ d46) + 32'hc4ac5665 + e0)) >> 32 - 23));
        
        //f = c ^ (b | (~d));
        //g = (7*i) % 16;
        b48 <= b47 + ((((a47 + (c47 ^ (b47 | (~d47))) + 32'hf4292244 + n47[63:32])) << 6) | (((a47 + (c47 ^ (b47 | (~d47))) + 32'hf4292244 + n47[63:32])) >> 32 - 6)); //g[0]
        b49 <= b48 + ((((a48 + (c48 ^ (b48 | (~d48))) + 32'h432aff97 + 0)) << 10) | (((a48 + (c48 ^ (b48 | (~d48))) + 32'h432aff97 + 0)) >> 32 - 10));
        b50 <= b49 + ((((a49 + (c49 ^ (b49 | (~d49))) + 32'hab9423a7 + e1)) << 15) | (((a49 + (c49 ^ (b49 | (~d49))) + 32'hab9423a7 + e1)) >> 32 - 15));
        b51 <= b50 + ((((a50 + (c50 ^ (b50 | (~d50))) + 32'hfc93a039 + 0)) << 21) | (((a50 + (c50 ^ (b50 | (~d50))) + 32'hfc93a039 + 0)) >> 32 - 21));
        
        b52 <= b51 + ((((a51 + (c51 ^ (b51 | (~d51))) + 32'h655b59c3 + 0)) << 6) | (((a51 + (c51 ^ (b51 | (~d51))) + 32'h655b59c3 + 0)) >> 32 - 6)); 
        b53 <= b52 + ((((a52 + (c52 ^ (b52 | (~d52))) + 32'h8f0ccc92 + 0)) << 10) | (((a52 + (c52 ^ (b52 | (~d52))) + 32'h8f0ccc92 + 0)) >> 32 - 10));
        b54 <= b53 + ((((a53 + (c53 ^ (b53 | (~d53))) + 32'hffeff47d + 0)) << 15) | (((a53 + (c53 ^ (b53 | (~d53))) + 32'hffeff47d + 0)) >> 32 - 15));
        b55 <= b54 + ((((a54 + (c54 ^ (b54 | (~d54))) + 32'h85845dd1 + n54[31:0])) << 21) | (((a54 + (c54 ^ (b54 | (~d54))) + 32'h85845dd1 + n54[31:0])) >> 32 - 21)); //g[1]
        
        b56 <= b55 + ((((a55 + (c55 ^ (b55 | (~d55))) + 32'h6fa87e4f + 0)) << 6) | (((a55 + (c55 ^ (b55 | (~d55))) + 32'h6fa87e4f + 0)) >> 32 - 6)); 
        b57 <= b56 + ((((a56 + (c56 ^ (b56 | (~d56))) + 32'hfe2ce6e0 + 0)) << 10) | (((a56 + (c56 ^ (b56 | (~d56))) + 32'hfe2ce6e0 + 0)) >> 32 - 10));
        b58 <= b57 + ((((a57 + (c57 ^ (b57 | (~d57))) + 32'ha3014314 + 0)) << 15) | (((a57 + (c57 ^ (b57 | (~d57))) + 32'ha3014314 + 0)) >> 32 - 15));
        b59 <= b58 + ((((a58 + (c58 ^ (b58 | (~d58))) + 32'h4e0811a1 + 0)) << 21) | (((a58 + (c58 ^ (b58 | (~d58))) + 32'h4e0811a1 + 0)) >> 32 - 21)); 
        
        b60 <= b59 + ((((a59 + (c59 ^ (b59 | (~d59))) + 32'hf7537e82 + 0)) << 6) | (((a59 + (c59 ^ (b59 | (~d59))) + 32'hf7537e82 + 0)) >> 32 - 6)); 
        b61 <= b60 + ((((a60 + (c60 ^ (b60 | (~d60))) + 32'hbd3af235 + 0)) << 10) | (((a60 + (c60 ^ (b60 | (~d60))) + 32'hbd3af235 + 0)) >> 32 - 10));
        b62 <= b61 + ((((a61 + (c61 ^ (b61 | (~d61))) + 32'h2ad7d2bb + e0)) << 15) | (((a61 + (c61 ^ (b61 | (~d61))) + 32'h2ad7d2bb + e0)) >> 32 - 15));
        b63 <= b62 + ((((a62 + (c62 ^ (b62 | (~d62))) + 32'heb86d391 + 0)) << 21) | (((a62 + (c62 ^ (b62 | (~d62))) + 32'heb86d391 + 0)) >> 32 - 21)); 
        
        a64 <= 32'h67452301 + a63;
        b64 <= 32'hefcdab89 + b63;
        c64 <= 32'h98badcfe + c63;
        d64 <= 32'h10325476 + d63;

end








endmodule
